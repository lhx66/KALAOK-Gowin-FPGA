parameter DIN_WIDTH = 16;
parameter COEFF_WIDTH = 12;
parameter DOUT_WIDTH = 16;
parameter NUM_CHN = 8;
parameter NUM_FACTOR = 1;
parameter TAPS_SIZE = 8;
parameter NUM_TDM = 1;
parameter COEFF_PATH = "./coeff.dat";
