`define MODULE_NAME Advanced_FIR_Filter_Top
`define fir_type_symmetry
