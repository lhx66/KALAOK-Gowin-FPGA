`define MODULE_NAME Equalizer_Ne
`define MUL_2;
