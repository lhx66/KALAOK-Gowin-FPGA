`define MODULE_NAME Equalizer_Po
`define MUL_2;
