`define MODULE_NAME Equalizer_Top
`define MUL_2;
