parameter BAND_SIZES = 10;
parameter GAIN_NUM = 5;
parameter COEFF_WIDTH = 16;
parameter DIN_WIDTH = 16;
parameter COEFFA_PATH = "./coeff_a.dat";
parameter COEFFB_PATH = "./coeff_b.dat";
